
module Verin (
	avalon_verin_0_conduit_end_clk_adc,
	avalon_verin_0_conduit_end_cs_n,
	avalon_verin_0_conduit_end_angle_barre,
	avalon_verin_0_conduit_end_pwm,
	avalon_verin_0_conduit_end_sens,
	clk_clk,
	reset_reset_n);	

	output		avalon_verin_0_conduit_end_clk_adc;
	output		avalon_verin_0_conduit_end_cs_n;
	input		avalon_verin_0_conduit_end_angle_barre;
	output		avalon_verin_0_conduit_end_pwm;
	output		avalon_verin_0_conduit_end_sens;
	input		clk_clk;
	input		reset_reset_n;
endmodule
